VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO oscilador
  CLASS BLOCK ;
  FOREIGN oscilador ;
  ORIGIN 47.020 -2.650 ;
  SIZE 37.060 BY 21.500 ;
  OBS
      LAYER nwell ;
        RECT -43.910 20.425 -36.170 22.030 ;
      LAYER pwell ;
        RECT -43.715 19.225 -36.365 20.135 ;
        RECT -43.570 19.035 -43.400 19.225 ;
      LAYER nwell ;
        RECT -43.850 16.735 -36.110 18.340 ;
        RECT -34.670 16.685 -30.150 18.290 ;
        RECT -28.740 16.565 -21.000 18.170 ;
        RECT -19.630 16.535 -13.730 18.140 ;
      LAYER pwell ;
        RECT -43.655 15.535 -36.305 16.445 ;
        RECT -43.510 15.345 -43.340 15.535 ;
        RECT -34.310 15.485 -30.440 16.395 ;
        RECT -34.310 15.465 -34.165 15.485 ;
        RECT -34.335 15.295 -34.165 15.465 ;
        RECT -28.545 15.365 -21.295 16.275 ;
        RECT -28.405 15.175 -28.235 15.365 ;
        RECT -19.435 15.335 -14.305 16.245 ;
        RECT -19.290 15.145 -19.120 15.335 ;
      LAYER nwell ;
        RECT -43.850 10.205 -36.110 11.810 ;
        RECT -34.520 10.285 -30.000 11.890 ;
        RECT -28.530 10.605 -20.790 12.210 ;
        RECT -19.110 10.715 -13.210 12.320 ;
      LAYER pwell ;
        RECT -43.655 9.005 -36.305 9.915 ;
        RECT -34.160 9.085 -30.290 9.995 ;
        RECT -28.335 9.405 -21.085 10.315 ;
        RECT -18.915 9.515 -13.785 10.425 ;
        RECT -28.195 9.215 -28.025 9.405 ;
        RECT -18.770 9.325 -18.600 9.515 ;
        RECT -34.160 9.065 -34.015 9.085 ;
        RECT -43.510 8.815 -43.340 9.005 ;
        RECT -34.185 8.895 -34.015 9.065 ;
      LAYER nwell ;
        RECT -43.770 6.235 -36.030 7.840 ;
      LAYER pwell ;
        RECT -43.575 5.035 -36.225 5.945 ;
        RECT -43.430 4.845 -43.260 5.035 ;
      LAYER li1 ;
        RECT -43.720 21.755 -36.360 21.925 ;
        RECT -43.630 20.615 -43.375 21.755 ;
        RECT -43.205 20.785 -42.875 21.585 ;
        RECT -42.705 20.955 -42.535 21.755 ;
        RECT -42.365 20.785 -42.035 21.585 ;
        RECT -41.865 20.955 -41.695 21.755 ;
        RECT -41.525 20.785 -41.195 21.585 ;
        RECT -41.025 20.955 -40.855 21.755 ;
        RECT -40.685 20.785 -40.355 21.585 ;
        RECT -40.185 20.955 -40.015 21.755 ;
        RECT -39.845 20.785 -39.515 21.585 ;
        RECT -39.345 20.955 -39.175 21.755 ;
        RECT -39.005 20.785 -38.675 21.585 ;
        RECT -38.505 20.955 -38.335 21.755 ;
        RECT -38.165 20.785 -37.835 21.585 ;
        RECT -37.665 20.955 -37.495 21.755 ;
        RECT -37.325 20.785 -36.995 21.585 ;
        RECT -43.205 20.585 -36.995 20.785 ;
        RECT -36.805 20.615 -36.450 21.755 ;
        RECT -43.210 20.195 -40.355 20.415 ;
        RECT -40.080 20.195 -39.600 20.585 ;
        RECT -38.120 20.580 -37.840 20.585 ;
        RECT -39.430 20.195 -37.415 20.395 ;
        RECT -39.845 20.025 -39.600 20.195 ;
        RECT -37.245 20.025 -36.995 20.585 ;
        RECT -43.630 19.855 -40.015 20.025 ;
        RECT -43.630 19.375 -43.295 19.855 ;
        RECT -43.125 19.205 -42.955 19.685 ;
        RECT -42.785 19.375 -42.455 19.855 ;
        RECT -42.285 19.205 -42.115 19.685 ;
        RECT -41.945 19.375 -41.615 19.855 ;
        RECT -41.445 19.205 -41.275 19.685 ;
        RECT -41.105 19.375 -40.775 19.855 ;
        RECT -40.605 19.205 -40.435 19.685 ;
        RECT -40.265 19.605 -40.015 19.855 ;
        RECT -39.845 19.775 -36.995 20.025 ;
        RECT -36.825 19.605 -36.450 20.025 ;
        RECT -40.265 19.375 -36.450 19.605 ;
        RECT -43.720 19.035 -36.360 19.205 ;
        RECT -43.660 18.065 -36.300 18.235 ;
        RECT -43.570 16.925 -43.315 18.065 ;
        RECT -43.145 17.095 -42.815 17.895 ;
        RECT -42.645 17.265 -42.475 18.065 ;
        RECT -42.305 17.095 -41.975 17.895 ;
        RECT -41.805 17.265 -41.635 18.065 ;
        RECT -41.465 17.095 -41.135 17.895 ;
        RECT -40.965 17.265 -40.795 18.065 ;
        RECT -40.625 17.095 -40.295 17.895 ;
        RECT -40.125 17.265 -39.955 18.065 ;
        RECT -39.785 17.095 -39.455 17.895 ;
        RECT -39.285 17.265 -39.115 18.065 ;
        RECT -38.945 17.095 -38.615 17.895 ;
        RECT -38.445 17.265 -38.275 18.065 ;
        RECT -38.105 17.095 -37.775 17.895 ;
        RECT -37.605 17.265 -37.435 18.065 ;
        RECT -37.265 17.095 -36.935 17.895 ;
        RECT -43.145 16.895 -36.935 17.095 ;
        RECT -36.745 16.925 -36.390 18.065 ;
        RECT -34.480 18.015 -30.340 18.185 ;
        RECT -34.225 17.215 -33.970 18.015 ;
        RECT -33.800 17.045 -33.470 17.845 ;
        RECT -33.300 17.215 -33.130 18.015 ;
        RECT -32.960 17.045 -32.630 17.845 ;
        RECT -32.460 17.215 -32.290 18.015 ;
        RECT -32.120 17.045 -31.790 17.845 ;
        RECT -31.620 17.215 -31.450 18.015 ;
        RECT -31.280 17.045 -30.950 17.845 ;
        RECT -30.780 17.215 -30.480 18.015 ;
        RECT -28.550 17.895 -21.190 18.065 ;
        RECT -43.150 16.505 -40.295 16.725 ;
        RECT -40.020 16.505 -39.540 16.895 ;
        RECT -39.370 16.505 -37.355 16.705 ;
        RECT -39.785 16.335 -39.540 16.505 ;
        RECT -37.185 16.335 -36.935 16.895 ;
        RECT -34.395 16.875 -30.425 17.045 ;
        RECT -43.570 16.165 -39.955 16.335 ;
        RECT -43.570 15.685 -43.235 16.165 ;
        RECT -43.065 15.515 -42.895 15.995 ;
        RECT -42.725 15.685 -42.395 16.165 ;
        RECT -42.225 15.515 -42.055 15.995 ;
        RECT -41.885 15.685 -41.555 16.165 ;
        RECT -41.385 15.515 -41.215 15.995 ;
        RECT -41.045 15.685 -40.715 16.165 ;
        RECT -40.545 15.515 -40.375 15.995 ;
        RECT -40.205 15.915 -39.955 16.165 ;
        RECT -39.785 16.085 -36.935 16.335 ;
        RECT -36.765 15.915 -36.390 16.335 ;
        RECT -34.395 16.285 -34.050 16.875 ;
        RECT -33.800 16.455 -30.945 16.705 ;
        RECT -30.745 16.285 -30.425 16.875 ;
        RECT -28.460 16.925 -28.145 17.725 ;
        RECT -27.975 17.095 -27.725 17.895 ;
        RECT -27.555 16.925 -27.305 17.725 ;
        RECT -27.135 17.095 -26.885 17.895 ;
        RECT -26.715 16.925 -26.465 17.725 ;
        RECT -26.295 17.095 -26.045 17.895 ;
        RECT -25.875 16.925 -25.625 17.725 ;
        RECT -25.455 17.095 -25.205 17.895 ;
        RECT -19.440 17.865 -13.920 18.035 ;
        RECT -25.035 17.555 -21.425 17.725 ;
        RECT -25.035 16.925 -24.785 17.555 ;
        RECT -28.460 16.715 -24.785 16.925 ;
        RECT -24.615 16.875 -24.365 17.385 ;
        RECT -24.195 17.045 -23.945 17.555 ;
        RECT -23.775 16.875 -23.525 17.385 ;
        RECT -23.355 17.045 -23.105 17.555 ;
        RECT -22.935 16.875 -22.685 17.385 ;
        RECT -22.515 17.045 -22.265 17.555 ;
        RECT -22.095 16.875 -21.845 17.385 ;
        RECT -21.675 17.045 -21.425 17.555 ;
        RECT -24.615 16.705 -21.275 16.875 ;
        RECT -28.190 16.335 -25.020 16.535 ;
        RECT -24.750 16.335 -22.010 16.535 ;
        RECT -34.395 16.095 -30.425 16.285 ;
        RECT -21.840 16.165 -21.275 16.705 ;
        RECT -19.345 16.845 -19.015 17.695 ;
        RECT -18.845 17.065 -18.675 17.865 ;
        RECT -18.505 16.845 -18.175 17.695 ;
        RECT -18.005 17.065 -17.835 17.865 ;
        RECT -17.585 16.845 -17.415 17.695 ;
        RECT -17.245 17.065 -16.915 17.865 ;
        RECT -16.745 16.845 -16.575 17.695 ;
        RECT -16.405 17.065 -16.075 17.865 ;
        RECT -15.905 16.845 -15.735 17.695 ;
        RECT -15.565 17.065 -15.235 17.865 ;
        RECT -15.065 16.845 -14.895 17.695 ;
        RECT -19.345 16.675 -17.845 16.845 ;
        RECT -17.585 16.675 -14.895 16.845 ;
        RECT -14.725 16.715 -14.395 17.865 ;
        RECT -19.300 16.305 -18.200 16.505 ;
        RECT -18.020 16.475 -17.845 16.675 ;
        RECT -18.020 16.305 -15.395 16.475 ;
        RECT -40.205 15.685 -36.390 15.915 ;
        RECT -43.660 15.345 -36.300 15.515 ;
        RECT -34.225 15.465 -33.970 15.925 ;
        RECT -33.800 15.635 -33.470 16.095 ;
        RECT -33.300 15.465 -33.130 15.925 ;
        RECT -32.960 15.635 -32.630 16.095 ;
        RECT -32.460 15.465 -32.290 15.925 ;
        RECT -32.120 15.635 -31.790 16.095 ;
        RECT -31.620 15.465 -31.450 15.925 ;
        RECT -31.280 15.635 -30.950 16.095 ;
        RECT -30.780 15.465 -30.475 15.925 ;
        RECT -34.480 15.295 -30.340 15.465 ;
        RECT -28.460 15.345 -28.185 16.165 ;
        RECT -28.015 15.985 -21.275 16.165 ;
        RECT -18.020 16.135 -17.845 16.305 ;
        RECT -15.150 16.135 -14.895 16.675 ;
        RECT -28.015 15.515 -27.685 15.985 ;
        RECT -27.515 15.345 -27.345 15.815 ;
        RECT -27.175 15.515 -26.845 15.985 ;
        RECT -26.675 15.345 -26.505 15.815 ;
        RECT -26.335 15.515 -26.005 15.985 ;
        RECT -25.835 15.345 -25.665 15.815 ;
        RECT -25.495 15.515 -25.165 15.985 ;
        RECT -24.995 15.345 -24.825 15.815 ;
        RECT -24.655 15.515 -24.325 15.985 ;
        RECT -24.155 15.345 -23.985 15.815 ;
        RECT -23.815 15.515 -23.485 15.985 ;
        RECT -23.315 15.345 -23.145 15.815 ;
        RECT -22.975 15.515 -22.645 15.985 ;
        RECT -22.475 15.345 -22.305 15.815 ;
        RECT -22.135 15.515 -21.805 15.985 ;
        RECT -19.265 15.965 -17.845 16.135 ;
        RECT -17.585 15.965 -14.895 16.135 ;
        RECT -21.635 15.345 -21.345 15.815 ;
        RECT -19.265 15.485 -19.095 15.965 ;
        RECT -28.550 15.175 -21.190 15.345 ;
        RECT -18.925 15.315 -18.595 15.795 ;
        RECT -18.425 15.490 -18.255 15.965 ;
        RECT -18.085 15.315 -17.755 15.795 ;
        RECT -17.585 15.485 -17.415 15.965 ;
        RECT -17.245 15.315 -16.915 15.795 ;
        RECT -16.745 15.485 -16.575 15.965 ;
        RECT -16.405 15.315 -16.075 15.795 ;
        RECT -15.905 15.485 -15.735 15.965 ;
        RECT -15.565 15.315 -15.235 15.795 ;
        RECT -15.065 15.485 -14.895 15.965 ;
        RECT -14.725 15.315 -14.395 16.115 ;
        RECT -19.440 15.145 -13.920 15.315 ;
        RECT -28.340 11.935 -20.980 12.105 ;
        RECT -18.920 12.045 -13.400 12.215 ;
        RECT -43.660 11.535 -36.300 11.705 ;
        RECT -34.330 11.615 -30.190 11.785 ;
        RECT -43.570 10.395 -43.315 11.535 ;
        RECT -43.145 10.565 -42.815 11.365 ;
        RECT -42.645 10.735 -42.475 11.535 ;
        RECT -42.305 10.565 -41.975 11.365 ;
        RECT -41.805 10.735 -41.635 11.535 ;
        RECT -41.465 10.565 -41.135 11.365 ;
        RECT -40.965 10.735 -40.795 11.535 ;
        RECT -40.625 10.565 -40.295 11.365 ;
        RECT -40.125 10.735 -39.955 11.535 ;
        RECT -39.785 10.565 -39.455 11.365 ;
        RECT -39.285 10.735 -39.115 11.535 ;
        RECT -38.945 10.565 -38.615 11.365 ;
        RECT -38.445 10.735 -38.275 11.535 ;
        RECT -38.105 10.565 -37.775 11.365 ;
        RECT -37.605 10.735 -37.435 11.535 ;
        RECT -37.265 10.565 -36.935 11.365 ;
        RECT -43.145 10.365 -36.935 10.565 ;
        RECT -36.745 10.395 -36.390 11.535 ;
        RECT -34.075 10.815 -33.820 11.615 ;
        RECT -33.650 10.645 -33.320 11.445 ;
        RECT -33.150 10.815 -32.980 11.615 ;
        RECT -32.810 10.645 -32.480 11.445 ;
        RECT -32.310 10.815 -32.140 11.615 ;
        RECT -31.970 10.645 -31.640 11.445 ;
        RECT -31.470 10.815 -31.300 11.615 ;
        RECT -31.130 10.645 -30.800 11.445 ;
        RECT -30.630 10.815 -30.330 11.615 ;
        RECT -28.250 10.965 -27.935 11.765 ;
        RECT -27.765 11.135 -27.515 11.935 ;
        RECT -27.345 10.965 -27.095 11.765 ;
        RECT -26.925 11.135 -26.675 11.935 ;
        RECT -26.505 10.965 -26.255 11.765 ;
        RECT -26.085 11.135 -25.835 11.935 ;
        RECT -25.665 10.965 -25.415 11.765 ;
        RECT -25.245 11.135 -24.995 11.935 ;
        RECT -24.825 11.595 -21.215 11.765 ;
        RECT -24.825 10.965 -24.575 11.595 ;
        RECT -28.250 10.755 -24.575 10.965 ;
        RECT -24.405 10.915 -24.155 11.425 ;
        RECT -23.985 11.085 -23.735 11.595 ;
        RECT -23.565 10.915 -23.315 11.425 ;
        RECT -23.145 11.085 -22.895 11.595 ;
        RECT -22.725 10.915 -22.475 11.425 ;
        RECT -22.305 11.085 -22.055 11.595 ;
        RECT -21.885 10.915 -21.635 11.425 ;
        RECT -21.465 11.085 -21.215 11.595 ;
        RECT -18.825 11.025 -18.495 11.875 ;
        RECT -18.325 11.245 -18.155 12.045 ;
        RECT -17.985 11.025 -17.655 11.875 ;
        RECT -17.485 11.245 -17.315 12.045 ;
        RECT -17.065 11.025 -16.895 11.875 ;
        RECT -16.725 11.245 -16.395 12.045 ;
        RECT -16.225 11.025 -16.055 11.875 ;
        RECT -15.885 11.245 -15.555 12.045 ;
        RECT -15.385 11.025 -15.215 11.875 ;
        RECT -15.045 11.245 -14.715 12.045 ;
        RECT -14.545 11.025 -14.375 11.875 ;
        RECT -24.405 10.745 -21.065 10.915 ;
        RECT -18.825 10.855 -17.325 11.025 ;
        RECT -17.065 10.855 -14.375 11.025 ;
        RECT -14.205 10.895 -13.875 12.045 ;
        RECT -34.245 10.475 -30.275 10.645 ;
        RECT -43.150 9.975 -40.295 10.195 ;
        RECT -40.020 9.975 -39.540 10.365 ;
        RECT -39.370 9.975 -37.355 10.175 ;
        RECT -39.785 9.805 -39.540 9.975 ;
        RECT -37.185 9.805 -36.935 10.365 ;
        RECT -34.245 9.885 -33.900 10.475 ;
        RECT -33.650 10.055 -30.795 10.305 ;
        RECT -30.595 9.885 -30.275 10.475 ;
        RECT -27.980 10.375 -24.810 10.575 ;
        RECT -24.540 10.375 -21.800 10.575 ;
        RECT -21.630 10.205 -21.065 10.745 ;
        RECT -18.780 10.485 -17.680 10.685 ;
        RECT -17.500 10.655 -17.325 10.855 ;
        RECT -17.500 10.485 -14.875 10.655 ;
        RECT -17.500 10.315 -17.325 10.485 ;
        RECT -14.630 10.315 -14.375 10.855 ;
        RECT -43.570 9.635 -39.955 9.805 ;
        RECT -43.570 9.155 -43.235 9.635 ;
        RECT -43.065 8.985 -42.895 9.465 ;
        RECT -42.725 9.155 -42.395 9.635 ;
        RECT -42.225 8.985 -42.055 9.465 ;
        RECT -41.885 9.155 -41.555 9.635 ;
        RECT -41.385 8.985 -41.215 9.465 ;
        RECT -41.045 9.155 -40.715 9.635 ;
        RECT -40.545 8.985 -40.375 9.465 ;
        RECT -40.205 9.385 -39.955 9.635 ;
        RECT -39.785 9.555 -36.935 9.805 ;
        RECT -36.765 9.385 -36.390 9.805 ;
        RECT -34.245 9.695 -30.275 9.885 ;
        RECT -40.205 9.155 -36.390 9.385 ;
        RECT -34.075 9.065 -33.820 9.525 ;
        RECT -33.650 9.235 -33.320 9.695 ;
        RECT -33.150 9.065 -32.980 9.525 ;
        RECT -32.810 9.235 -32.480 9.695 ;
        RECT -32.310 9.065 -32.140 9.525 ;
        RECT -31.970 9.235 -31.640 9.695 ;
        RECT -31.470 9.065 -31.300 9.525 ;
        RECT -31.130 9.235 -30.800 9.695 ;
        RECT -30.630 9.065 -30.325 9.525 ;
        RECT -28.250 9.385 -27.975 10.205 ;
        RECT -27.805 10.025 -21.065 10.205 ;
        RECT -18.745 10.145 -17.325 10.315 ;
        RECT -17.065 10.145 -14.375 10.315 ;
        RECT -27.805 9.555 -27.475 10.025 ;
        RECT -27.305 9.385 -27.135 9.855 ;
        RECT -26.965 9.555 -26.635 10.025 ;
        RECT -26.465 9.385 -26.295 9.855 ;
        RECT -26.125 9.555 -25.795 10.025 ;
        RECT -25.625 9.385 -25.455 9.855 ;
        RECT -25.285 9.555 -24.955 10.025 ;
        RECT -24.785 9.385 -24.615 9.855 ;
        RECT -24.445 9.555 -24.115 10.025 ;
        RECT -23.945 9.385 -23.775 9.855 ;
        RECT -23.605 9.555 -23.275 10.025 ;
        RECT -23.105 9.385 -22.935 9.855 ;
        RECT -22.765 9.555 -22.435 10.025 ;
        RECT -22.265 9.385 -22.095 9.855 ;
        RECT -21.925 9.555 -21.595 10.025 ;
        RECT -21.425 9.385 -21.135 9.855 ;
        RECT -18.745 9.665 -18.575 10.145 ;
        RECT -18.405 9.495 -18.075 9.975 ;
        RECT -17.905 9.670 -17.735 10.145 ;
        RECT -17.565 9.495 -17.235 9.975 ;
        RECT -17.065 9.665 -16.895 10.145 ;
        RECT -16.725 9.495 -16.395 9.975 ;
        RECT -16.225 9.665 -16.055 10.145 ;
        RECT -15.885 9.495 -15.555 9.975 ;
        RECT -15.385 9.665 -15.215 10.145 ;
        RECT -15.045 9.495 -14.715 9.975 ;
        RECT -14.545 9.665 -14.375 10.145 ;
        RECT -14.205 9.495 -13.875 10.295 ;
        RECT -28.340 9.215 -20.980 9.385 ;
        RECT -18.920 9.325 -13.400 9.495 ;
        RECT -43.660 8.815 -36.300 8.985 ;
        RECT -34.330 8.895 -30.190 9.065 ;
        RECT -43.580 7.565 -36.220 7.735 ;
        RECT -43.490 6.425 -43.235 7.565 ;
        RECT -43.065 6.595 -42.735 7.395 ;
        RECT -42.565 6.765 -42.395 7.565 ;
        RECT -42.225 6.595 -41.895 7.395 ;
        RECT -41.725 6.765 -41.555 7.565 ;
        RECT -41.385 6.595 -41.055 7.395 ;
        RECT -40.885 6.765 -40.715 7.565 ;
        RECT -40.545 6.595 -40.215 7.395 ;
        RECT -40.045 6.765 -39.875 7.565 ;
        RECT -39.705 6.595 -39.375 7.395 ;
        RECT -39.205 6.765 -39.035 7.565 ;
        RECT -38.865 6.595 -38.535 7.395 ;
        RECT -38.365 6.765 -38.195 7.565 ;
        RECT -38.025 6.595 -37.695 7.395 ;
        RECT -37.525 6.765 -37.355 7.565 ;
        RECT -37.185 6.595 -36.855 7.395 ;
        RECT -43.065 6.395 -36.855 6.595 ;
        RECT -36.665 6.425 -36.310 7.565 ;
        RECT -43.070 6.005 -40.215 6.225 ;
        RECT -39.940 6.005 -39.460 6.395 ;
        RECT -39.290 6.005 -37.275 6.205 ;
        RECT -39.705 5.835 -39.460 6.005 ;
        RECT -37.105 5.835 -36.855 6.395 ;
        RECT -43.490 5.665 -39.875 5.835 ;
        RECT -43.490 5.185 -43.155 5.665 ;
        RECT -42.985 5.015 -42.815 5.495 ;
        RECT -42.645 5.185 -42.315 5.665 ;
        RECT -42.145 5.015 -41.975 5.495 ;
        RECT -41.805 5.185 -41.475 5.665 ;
        RECT -41.305 5.015 -41.135 5.495 ;
        RECT -40.965 5.185 -40.635 5.665 ;
        RECT -40.465 5.015 -40.295 5.495 ;
        RECT -40.125 5.415 -39.875 5.665 ;
        RECT -39.705 5.585 -36.855 5.835 ;
        RECT -36.685 5.415 -36.310 5.835 ;
        RECT -40.125 5.185 -36.310 5.415 ;
        RECT -43.580 4.845 -36.220 5.015 ;
      LAYER met1 ;
        RECT -44.960 24.140 -24.470 24.150 ;
        RECT -44.960 24.130 -20.670 24.140 ;
        RECT -44.960 23.630 -20.350 24.130 ;
        RECT -44.960 22.980 -44.520 23.630 ;
        RECT -24.480 23.620 -20.350 23.630 ;
        RECT -20.750 23.600 -20.350 23.620 ;
        RECT -44.960 22.450 -44.510 22.980 ;
        RECT -44.950 20.430 -44.510 22.450 ;
        RECT -43.720 21.950 -36.360 22.080 ;
        RECT -43.720 21.710 -33.820 21.950 ;
        RECT -43.720 21.600 -36.360 21.710 ;
        RECT -39.350 20.580 -35.550 20.720 ;
        RECT -47.020 20.380 -42.880 20.430 ;
        RECT -39.350 20.390 -39.180 20.580 ;
        RECT -35.800 20.390 -35.550 20.580 ;
        RECT -47.020 20.190 -40.430 20.380 ;
        RECT -39.900 20.290 -35.550 20.390 ;
        RECT -39.900 20.190 -35.540 20.290 ;
        RECT -44.950 16.720 -44.510 20.190 ;
        RECT -43.210 20.140 -40.430 20.190 ;
        RECT -43.720 18.880 -36.360 19.360 ;
        RECT -43.660 18.260 -36.300 18.390 ;
        RECT -35.860 18.260 -35.540 20.190 ;
        RECT -34.510 18.340 -34.160 21.710 ;
        RECT -20.750 20.205 -20.370 23.600 ;
        RECT -20.750 20.200 -20.365 20.205 ;
        RECT -20.800 19.820 -20.320 20.200 ;
        RECT -34.510 18.260 -30.340 18.340 ;
        RECT -43.660 18.150 -30.340 18.260 ;
        RECT -28.550 18.150 -21.190 18.220 ;
        RECT -43.660 17.920 -21.190 18.150 ;
        RECT -43.660 17.910 -30.340 17.920 ;
        RECT -36.620 17.890 -30.340 17.910 ;
        RECT -35.860 16.730 -35.540 17.890 ;
        RECT -34.480 17.860 -30.340 17.890 ;
        RECT -28.550 17.740 -21.190 17.920 ;
        RECT -20.750 17.670 -20.365 19.820 ;
        RECT -19.440 17.710 -13.920 18.190 ;
        RECT -44.950 16.700 -42.860 16.720 ;
        RECT -35.890 16.700 -35.510 16.730 ;
        RECT -44.950 16.680 -41.980 16.700 ;
        RECT -39.850 16.690 -33.570 16.700 ;
        RECT -41.730 16.680 -33.570 16.690 ;
        RECT -44.950 16.530 -33.570 16.680 ;
        RECT -20.745 16.650 -20.365 17.670 ;
        RECT -30.460 16.540 -27.940 16.630 ;
        RECT -44.950 16.520 -44.510 16.530 ;
        RECT -43.980 16.510 -33.570 16.530 ;
        RECT -42.980 16.500 -33.570 16.510 ;
        RECT -42.980 16.490 -40.980 16.500 ;
        RECT -43.660 15.530 -36.300 15.670 ;
        RECT -35.860 15.530 -35.540 16.500 ;
        RECT -30.650 16.400 -27.940 16.540 ;
        RECT -20.750 16.500 -20.360 16.650 ;
        RECT -12.670 16.510 -10.140 16.520 ;
        RECT -21.390 16.300 -18.230 16.500 ;
        RECT -15.140 16.060 -10.140 16.510 ;
        RECT -15.140 16.050 -12.610 16.060 ;
        RECT -34.480 15.530 -30.340 15.620 ;
        RECT -43.660 15.480 -30.340 15.530 ;
        RECT -28.550 15.480 -21.190 15.500 ;
        RECT -43.660 15.420 -21.190 15.480 ;
        RECT -19.440 15.420 -13.920 15.470 ;
        RECT -43.660 15.300 -13.920 15.420 ;
        RECT -43.660 15.190 -36.300 15.300 ;
        RECT -41.480 12.890 -41.250 14.390 ;
        RECT -41.480 12.710 -39.610 12.890 ;
        RECT -39.830 11.860 -39.650 12.710 ;
        RECT -43.660 11.700 -36.300 11.860 ;
        RECT -35.860 11.700 -35.540 15.300 ;
        RECT -34.480 15.260 -13.920 15.300 ;
        RECT -34.480 15.140 -30.340 15.260 ;
        RECT -28.550 15.100 -13.920 15.260 ;
        RECT -28.550 15.020 -21.190 15.100 ;
        RECT -19.440 14.990 -13.920 15.100 ;
        RECT -28.340 12.130 -20.980 12.260 ;
        RECT -18.920 12.130 -13.400 12.370 ;
        RECT -28.340 12.040 -13.400 12.130 ;
        RECT -30.350 11.940 -13.400 12.040 ;
        RECT -34.330 11.900 -13.400 11.940 ;
        RECT -34.330 11.780 -20.980 11.900 ;
        RECT -18.920 11.890 -13.400 11.900 ;
        RECT -34.330 11.770 -27.800 11.780 ;
        RECT -34.330 11.700 -30.190 11.770 ;
        RECT -43.660 11.520 -30.190 11.700 ;
        RECT -43.660 11.380 -36.300 11.520 ;
        RECT -44.240 10.190 -40.310 10.200 ;
        RECT -45.450 9.990 -40.310 10.190 ;
        RECT -39.830 10.020 -39.650 11.380 ;
        RECT -38.400 10.150 -37.960 10.160 ;
        RECT -35.860 10.150 -35.540 11.520 ;
        RECT -34.330 11.460 -30.190 11.520 ;
        RECT -14.630 10.670 -12.140 10.680 ;
        RECT -30.625 10.270 -30.245 10.330 ;
        RECT -29.410 10.270 -21.800 10.560 ;
        RECT -20.070 10.490 -18.450 10.640 ;
        RECT -21.170 10.480 -18.450 10.490 ;
        RECT -21.170 10.330 -19.550 10.480 ;
        RECT -14.630 10.310 -9.960 10.670 ;
        RECT -12.450 10.300 -9.960 10.310 ;
        RECT -30.625 10.240 -21.800 10.270 ;
        RECT -35.190 10.150 -33.410 10.210 ;
        RECT -38.400 10.060 -33.410 10.150 ;
        RECT -38.400 10.010 -34.490 10.060 ;
        RECT -38.000 10.000 -34.490 10.010 ;
        RECT -45.450 9.980 -42.600 9.990 ;
        RECT -45.450 9.310 -45.020 9.980 ;
        RECT -30.625 9.950 -29.090 10.240 ;
        RECT -30.625 9.890 -30.245 9.950 ;
        RECT -18.920 9.540 -13.400 9.650 ;
        RECT -45.460 9.080 -45.020 9.310 ;
        RECT -28.340 9.310 -13.400 9.540 ;
        RECT -28.340 9.290 -20.980 9.310 ;
        RECT -30.430 9.220 -20.980 9.290 ;
        RECT -45.460 7.680 -45.030 9.080 ;
        RECT -43.660 9.010 -36.300 9.140 ;
        RECT -34.330 9.060 -20.980 9.220 ;
        RECT -18.920 9.170 -13.400 9.310 ;
        RECT -34.330 9.020 -27.880 9.060 ;
        RECT -34.330 9.010 -30.190 9.020 ;
        RECT -43.660 8.740 -30.190 9.010 ;
        RECT -43.660 8.660 -36.300 8.740 ;
        RECT -45.470 6.930 -45.030 7.680 ;
        RECT -43.580 7.750 -36.220 7.890 ;
        RECT -43.580 7.430 -34.760 7.750 ;
        RECT -43.580 7.410 -36.220 7.430 ;
        RECT -45.470 6.230 -45.040 6.930 ;
        RECT -45.470 6.220 -40.210 6.230 ;
        RECT -46.240 6.010 -40.210 6.220 ;
        RECT -39.830 6.220 -39.470 6.240 ;
        RECT -39.830 6.210 -39.290 6.220 ;
        RECT -38.870 6.210 -35.250 6.230 ;
        RECT -46.240 5.990 -45.040 6.010 ;
        RECT -39.830 6.000 -35.250 6.210 ;
        RECT -45.470 3.140 -45.040 5.990 ;
        RECT -39.490 5.980 -35.250 6.000 ;
        RECT -39.130 5.970 -35.250 5.980 ;
        RECT -38.830 5.170 -38.560 5.970 ;
        RECT -43.580 4.690 -36.220 5.170 ;
        RECT -38.810 4.530 -38.540 4.690 ;
        RECT -38.810 4.520 -35.970 4.530 ;
        RECT -35.750 4.520 -35.250 5.970 ;
        RECT -38.810 4.190 -35.230 4.520 ;
        RECT -36.200 4.180 -35.230 4.190 ;
        RECT -45.470 3.130 -24.580 3.140 ;
        RECT -45.470 3.110 -22.380 3.130 ;
        RECT -45.470 2.680 -19.560 3.110 ;
        RECT -24.680 2.670 -19.560 2.680 ;
        RECT -22.490 2.650 -19.560 2.670 ;
      LAYER met2 ;
        RECT -20.750 19.770 -20.370 20.250 ;
        RECT -36.550 19.210 -35.060 19.230 ;
        RECT -36.550 18.970 -35.020 19.210 ;
        RECT -43.140 16.700 -40.350 16.730 ;
        RECT -44.770 16.690 -40.350 16.700 ;
        RECT -44.790 16.530 -40.350 16.690 ;
        RECT -44.790 16.500 -41.980 16.530 ;
        RECT -44.790 14.390 -44.400 16.500 ;
        RECT -44.790 14.210 -41.290 14.390 ;
        RECT -39.840 13.240 -39.620 16.670 ;
        RECT -45.020 13.220 -43.620 13.230 ;
        RECT -45.020 13.210 -42.260 13.220 ;
        RECT -41.220 13.210 -39.590 13.240 ;
        RECT -45.020 13.090 -39.590 13.210 ;
        RECT -45.010 13.070 -40.960 13.090 ;
        RECT -39.840 13.080 -39.620 13.090 ;
        RECT -45.010 12.340 -44.570 13.070 ;
        RECT -42.360 13.060 -40.960 13.070 ;
        RECT -45.010 12.020 -44.560 12.340 ;
        RECT -45.000 10.200 -44.560 12.020 ;
        RECT -45.000 10.180 -44.500 10.200 ;
        RECT -45.000 10.150 -42.580 10.180 ;
        RECT -40.400 10.160 -37.390 10.180 ;
        RECT -41.570 10.150 -37.390 10.160 ;
        RECT -45.000 10.010 -37.390 10.150 ;
        RECT -44.750 10.000 -37.390 10.010 ;
        RECT -43.190 9.980 -39.580 10.000 ;
        RECT -43.190 9.970 -41.200 9.980 ;
        RECT -35.860 5.980 -35.540 16.730 ;
        RECT -35.270 15.460 -35.020 18.970 ;
        RECT -21.580 17.710 -19.240 18.140 ;
        RECT -22.840 16.530 -20.440 16.540 ;
        RECT -24.760 16.350 -20.440 16.530 ;
        RECT -24.760 16.340 -20.350 16.350 ;
        RECT -24.760 16.330 -22.040 16.340 ;
        RECT -35.270 15.230 -34.140 15.460 ;
        RECT -20.720 14.340 -20.350 16.340 ;
        RECT -29.610 12.870 -24.830 12.900 ;
        RECT -29.610 12.680 -20.940 12.870 ;
        RECT -35.270 11.580 -34.250 11.740 ;
        RECT -35.270 7.480 -34.830 11.580 ;
        RECT -29.600 10.560 -29.370 12.680 ;
        RECT -25.720 12.650 -20.940 12.680 ;
        RECT -21.210 12.640 -20.970 12.650 ;
        RECT -29.600 10.550 -26.590 10.560 ;
        RECT -29.600 10.380 -24.860 10.550 ;
        RECT -27.850 10.370 -24.860 10.380 ;
        RECT -21.300 10.490 -21.110 10.910 ;
        RECT -20.680 10.490 -20.450 14.340 ;
        RECT -21.300 10.440 -20.450 10.490 ;
        RECT -21.300 10.330 -20.460 10.440 ;
        RECT -20.070 9.440 -19.550 10.420 ;
        RECT -34.320 5.020 -33.960 9.100 ;
        RECT -20.080 8.560 -19.550 9.440 ;
        RECT -20.090 8.310 -19.550 8.560 ;
        RECT -20.090 6.780 -19.560 8.310 ;
        RECT -36.640 4.750 -33.960 5.020 ;
        RECT -34.320 4.740 -33.960 4.750 ;
        RECT -20.110 6.650 -19.560 6.780 ;
        RECT -20.110 3.040 -19.580 6.650 ;
      LAYER met3 ;
        RECT -21.210 16.500 -20.910 16.610 ;
        RECT -21.210 16.300 -20.900 16.500 ;
        RECT -21.200 12.950 -20.900 16.300 ;
        RECT -21.200 12.640 -20.870 12.950 ;
  END
END oscilador
END LIBRARY

